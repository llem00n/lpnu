LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TSG IS
  PORT (
    RST : OUT STD_LOGIC;
    PUSK : OUT STD_LOGIC;
    X : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    CLK : OUT STD_LOGIC
  );
END TSG;
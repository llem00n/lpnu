LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ARCHITECTURE Implementation OF TSG IS
BEGIN
  PROCESS
  BEGIN
    WAIT;
  END PROCESS;
END Implementation;